-- Laboratório 07 -> Função principal.
Library IEEE;
use ieee.std_logic_1164.all;

entity Lab07 is
    port (

    );
end Lab07;


architecture struct of Lab07 is

--signals 

--components

    begin 



    end struct;
