-- Laboratório 05 -> Função principal.
Library IEEE;
use ieee.std_logic_1164.all;

entity Lab05 is
    port (
      
    );
end Lab05;