-- Função principal do Laboratório 03.
-- Laboratório 03 -> Função principal.
Library IEEE;
use ieee.std_logic_1164.all;

entity Lab03 is
    port (
        pb0: in std_logic;
        pb1: in std_logic;
        sw: in std_logic_vector (7 downto 0);
        leds: out std_logic_vector (7 downto 0);
        hex0: out std_logic_vector (3 downto 0);
        hex1: out std_logic_vector (3 downto 0)
    );
end Lab03;

architecture struct of Lab03 is
    begin 
        

    end struct;