-- Projete e implemente um conversor PISO (Parallel-in, Serial-out) de 8 bits.
