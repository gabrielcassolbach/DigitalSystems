-- Projete e implemente um conversor PISO (Serial-in, Parallel-out) de 8 bits.
