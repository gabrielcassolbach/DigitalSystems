--Função principal do laboratório 02.
Library IEEE;
use ieee.std_logic_1164.all;


entity Lab02_1 is 
	port (
		
	);
end Lab02_1;


--passo 1: gerar o deslocamento de bits utilizando um registrador paralelo
-- precisa-se de: 4 flip-flops-d, 

architecture struct of Lab02_1 is
    begin

    end struct;